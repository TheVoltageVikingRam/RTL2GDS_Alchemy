`ifndef SANDPIPER_GEN_VH
`define SANDPIPER_GEN_VH

// Clock and reset signals
`define BOGUS_USE(var)

`endif
