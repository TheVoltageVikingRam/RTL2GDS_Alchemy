module dff_asyncres_syncres (input clk, input async_reset, input sync_res, input d, output reg q);
always @ (posedge clk, posedge async_reset)
begin
	if (async_reset)
		q<=1'b0;
	else if (sync_reset)
		q<=1'b0;
	else
		q<=d;
end
endmodule
