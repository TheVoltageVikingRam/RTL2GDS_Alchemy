***MODEL Descriptions***
***NETLIST Description***

M1 out in vdd vdd pmos W=0.375u L=0.25u
M2 our in 0 0 nmos W=0.375u L=0.25u

cload out 0 10f

Vdd vdd 0 2.5
Vin in 0 2.5

***SIMULATION Commands***


.op
.dc vin 0 2.5 0.05
*** .include tsmc_025um_model.mod ***
.LIB "tsmc_025um_model.mod" CMOS_MODELS

.end
