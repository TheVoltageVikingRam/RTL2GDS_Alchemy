`ifndef SP_VERILOG_VH
`define SP_VERILOG_VH
`endif
